module registerFile();

endmodule
